** sch_path:
*+ /home/grigorii/projects/OpenLane/pdks/sky130A/libs.tech/xschem/sky130_tests/test_vpp_cap.sch
**.subckt test_vpp_cap
I1 0 G pwl 0 0 1000n 0 1010n 100n
R1 G REF 1G m=1
I3 0 G2 pwl 0 0 1000n 0 1010n 100n
R3 G2 REF 1G m=1
C1 G2 0 0.148p m=1
V1 REF 0 -2
XC2 G 0 0 0 sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3m4_shieldm5 W=1 L=1 mult=1 m=1
**** begin user architecture code


.control
tran 10n 6u
**** plot g g2
**** write test_vpp_cap.raw
hardcopy test_vpp_cap.svg g g2
.endc



** opencircuitdesign pdks install
.lib /home/grigorii/projects/OpenLane/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
**.ends
.end
