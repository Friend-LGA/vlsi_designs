** sch_path:
*+ /home/grigorii_lutkov/Projects/OpenLane/pdks/sky130A/libs.tech/xschem/sky130_tests/test_bipolar.sch
**.subckt test_bipolar
XQ1 net2 net1 E1 sky130_fd_pr__pnp_05v5_W3p40L3p40
Vc1 net2 0 0
.save  i(vc1)
Vb1 net1 0 0
.save  i(vb1)
I0 0 net3 0
Ve1 net3 E1 0
.save  i(ve1)
**** begin user architecture code


.control
save all
dc i0 5n 5u 0.05u
* tran 1n 2u
****plot vc1#branch / vb1#branch
****plot e1
hardcopy test_bipolar.svg vc1#branch / vb1#branch
.endc



** opencircuitdesign pdks install
.lib /home/grigorii_lutkov/Projects/OpenLane/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt

**** end user architecture code
**.ends
.end
