** sch_path:
*+ /home/grigorii_lutkov/Projects/OpenLane/pdks/sky130A/libs.tech/xschem/sky130_tests/test_varactor.sch
**.subckt test_varactor
I1 0 G pwl 0 0 1n 100n
R1 G REF 1G m=1
I2 0 G1 pwl 0 0 1n 100n
R2 G1 REF 1G m=1
I3 0 G2 pwl 0 0 1n 100n
R3 G2 REF 1G m=1
C1 G2 0 0.19p m=1
V1 REF 0 -2
XM1 0 G1 0 0 sky130_fd_pr__nfet_01v8_lvt L=5 W=5 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)'
+ ps='2 * (W + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
I4 0 G3 pwl 0 0 1n 100n
R4 G3 REF 1G m=1
C2 G3 0 q='v(g3) * 0.19p' m=1
XC4 G 0 0 sky130_fd_pr__cap_var_lvt W=5 L=5 VM=1 m=1
**** begin user architecture code


.control
tran 10n 9u
****plot g g1 g2 g3
****plot '100n/deriv(g)' vs v(g) ylimit 0 0.3p
****plot '100n/deriv(g1)' vs v(g1) ylimit 0 0.3p
****write test_varactor.raw
hardcopy test_varactor.svg g g1 g2 g3
.endc



** opencircuitdesign pdks install
.lib /home/grigorii_lutkov/Projects/OpenLane/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
**.ends
.end
